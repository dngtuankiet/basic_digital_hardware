/*
Date: 11/05/2019
Name: Dang Tuan Kiet
Description: 4-bit Carray Look Ahead Adder
*/

module CLA_4bit(i_a,
					      i_b,
				      	 i_ci,
				      	 o_s,
				      	 o_co
					      );

input [3:0] i_a;
input [3:0] i_b;
input i_ci;
output [3:0] o_s;
output o_co;

wire [8:0] s1;
wire [18:0] s2;
wire [8:0] s3;

//S1
assign
s1[8] = ~i_ci,
s1[7] = ~(i_a[0] | i_b[0]),
s1[6] = ~(i_a[0] & i_b[0]),

s1[5] = ~(i_a[1] | i_b[1]),
s1[4] = ~(i_a[1] & i_b[1]),

s1[3] = ~(i_a[2] | i_b[2]),
s1[2] = ~(i_a[2] & i_b[2]),

s1[1] = ~(i_a[3] | i_b[3]),
s1[0] = ~(i_a[3] & i_b[3]);

//S2
assign
s2[18] = ~s1[8],
s2[17] = ~s1[7] & s1[6],

s2[16] = s1[8] & s1[6],
s2[15] = s1[7],

s2[14] = ~s1[5] & s1[4],
s2[13] = ((s1[8] & s1[6]) & s1[4]),
s2[12] = s1[4] & s1[7],
s2[11] = s1[5],

s2[10] = ~s1[3] & s1[2],
s2[9]  = ((s1[8] & s1[6]) & (s1[4] & s1[2])),
s2[8]  = s1[4] & s1[2] & s1[7],
s2[7] = s1[2] & s1[5],
s2[6] = s1[3],

s2[5] = ~s1[1] & s1[0],
s2[4] = (((s1[8] & s1[6]) & s1[4]) & s1[2]) & s1[0],
s2[3] = ((s1[4] & s1[2]) & s1[0]) & s1[7],
s2[2] = (s1[2] & s1[0]) & s1[5],
s2[1] = s1[0] & s1[3],
s2[0] = s1[1];

//S3
assign
s3[8] = s2[18],
s3[7] = s2[17],

s3[6] = ~(s2[16] | s2[15]),
s3[5] = s2[14],

s3[4] = ~((s2[13] | s2[12]) | s2[11]),
s3[3] = s2[10],

s3[2] = ~(((s2[9] | s2[8]) | s2[7]) | s2[6]),
s3[1] = s2[5],

s3[0] = ~((s2[4] | s2[3]) | ((s2[2] | s2[1]) | s2[0]));

//Output
assign
o_s[0] = s3[8] ^ s3[7],
o_s[1] = s3[6] ^ s3[5],
o_s[2] = s3[4] ^ s3[3],
o_s[3] = s3[2] ^ s3[1],
o_co = s3[0];

endmodule
